`timescale 10ns/1ns
module fsub_TB;
reg ain,bin,cin; //???????
wire sum,borrow; //?????????
initial //?????????? initial ??
    begin //initial ????????? begin end
        ain=0;bin=0;cin=0; //??????? T=0 ????a,b,c ???? 0??????
        #10 ain=0;bin=0;cin=1; // T=100ns ?????????? 001
        #10 ain=0;bin=1;cin=0; // T=200ns ?????????? 010
        #10 ain=0;bin=1;cin=1; // T=300ns ?????????? 011
        #10 ain=1;bin=0;cin=0; // T=400ns ?????????? 100
        #10 ain=1;bin=0;cin=1; // T=500ns ?????????? 101
        #10 ain=1;bin=1;cin=0; // T=600ns ?????????? 110
        #10 ain=1;bin=1;cin=1; // T=700ns ?????????? 111
        #10 $stop; //?????????????,???? Stop ???????
    end
fsub m1(.SUM(sum),.BORROW(borrow),.A(ain),.B(bin),.C(cin)); //????

endmodule

