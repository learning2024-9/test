`timescale 10ns/1ns
module fsub_4b_TB;
reg [3:0]A,B; //4 ????
reg CIN; //?????
wire [3:0] SUM; //???
wire BORROW; //?????
initial //????
    begin
        A=4'b0000;B=4'b1100;CIN=0; //?????? 1?b1?B ???A ??
        #10 A=4'b0001; //A ?? 4?b0000-4?b1111
        #10 A=4'b0010; #10 A=4'b0011; #10 A=4'b0100; #10 A=4'b0101;
        #10 A=4'b0110; #10 A=4'b0111; #10 A=4'b1000; #10 A=4'b1001;
        #10 A=4'b1010; #10 A=4'b1011; #10 A=4'b1100; #10 A=4'b1101;
        #10 A=4'b1110; #10 A=4'b1111;
        //?????? 1?b1?A ???B ?? 4?b0000-4?b1111
        #10 A=4'b1100; B=4'b0000; CIN=1'b1;
        #10 B=4'b0001; #10 B=4'b0010; #10 B=4'b0011; #10 B=4'b0100;
        #10 B=4'b0101; #10 B=4'b0110; #10 B=4'b0111; #10 B=4'b1000;
        #10 B=4'b1001; #10 B=4'b1010; #10 B=4'b1011; #10 B=4'b1100;
        #10 B=4'b1101; #10 B=4'b1110; #10 B=4'b1111; 
        #10 $stop; //????
    end
fsub_4b m0(SUM,BORROW,A,B,CIN); //??????
endmodule